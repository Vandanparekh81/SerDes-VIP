//---------------------------------------------------------------------------------------------//
// File Name : serdes_same_data_for_tx_rx_sequence.sv
// Author Name : Vandan Parekh
// Propetier Name : ASICraft Technologies LLP.
// Decription : This is serdes_same_data_for_tx_rx_sequence in this sequence it generates same 
// data of Tx0 for Rx0_p for example if Tx0 generated data is 0001110001 then Rx0_p generated 
// data is 0001110001 
//---------------------------------------------------------------------------------------------//

class serdes_same_data_for_tx_rx_sequence extends serdes_base_sequence;

  // Factory registration of sequence class
  `uvm_object_utils(serdes_same_data_for_tx_rx_sequence);

  // Properties declaration of sequence class
  bit is_parallel; // Indicates if the sequence is for a parallel or serial agent
  event synchro_seq; // Event for synchronization between two sequence

  // Constructor of sequence class
  function new(string name = "serdes_same_data_for_tx_rx_sequence");
    super.new(name);
  endfunction : new

  // Pre body task
  virtual task pre_body();
    super.pre_body();
  endtask : pre_body

  // This body task generate transactions and send to arbitration of sequencer and this task also differentiate between generate serial transaction and parallel transaction
  virtual task body();
    req = serdes_transaction::type_id::create("req"); // Creation of transaction packet
    // IF is_parallel is 1 then it will generate parallel data otherwise it will generate serial data
    if(is_parallel) begin
        `uvm_info("BODY", $sformatf("Begin of parallel"), UVM_LOW)
      // For parallel agent: Generate one transaction with randomized Tx0
      repeat(parallel_transaction_count) begin
        `uvm_info("BODY", $sformatf("Begin of parallel  2"), UVM_LOW)
        start_item(req);
        `uvm_info("BODY", $sformatf("Begin of parallel 3"), UVM_LOW)
        assert(req.randomize() with { Tx0 != 0; });// Ensure non-zero for testing
        uvm_config_db#(int)::set(null, "*", "same_data", req.Tx0);
        -> synchro_seq;
        `uvm_info("BODY", $sformatf("Parallel transaction: Tx0 in Binary=%b | Tx0 in Decimal = %0d", req.Tx0,req.Tx0), UVM_LOW)
        finish_item(req); // This task will return if driver provide item_done
        `uvm_info("BODY", $sformatf("AFTER Finish Item Parallel transaction: Tx0 in Binary=%b | Tx0 in Decimal = %0d", req.Tx0,req.Tx0), UVM_LOW)
      end
    end

    // If is_parallel is 0 means i have to generate serial transactions 
    else begin
        `uvm_info("BODY", $sformatf("Begin of Serial"), UVM_LOW)
      // For serial agent: Generate 1 transactions for Rx0_p and Rx0_n
      repeat(serial_transaction_count) begin // WIDTH=10 for serial bits
        `uvm_info("BODY", $sformatf("Begin of Serial 2"), UVM_LOW)
        start_item(req); 
        `uvm_info("BODY", $sformatf("Begin of Serial 3"), UVM_LOW)
        @(synchro_seq);
        if(!uvm_config_db#(int)::get(null, "*", "same_data", req.Rx0_p))
          `uvm_fatal("NO_SAMEDATA",{"Same data should be set for sequence 1: ",get_full_name()});
        //assert(req.randomize() with { Rx0_p != 0; }); // Equal distribution for 0 and 1
        `uvm_info("BODY", $sformatf("Serial transaction: Rx0_p=%b (%0d)",req.Rx0_p, req.Rx0_p), UVM_LOW)
        finish_item(req); // This task will return if driver provide item_done
        `uvm_info("BODY", $sformatf("After Finish item Serial transaction: Rx0_p=%b (%0d)",req.Rx0_p, req.Rx0_p), UVM_LOW)
      end
    end
        `uvm_info("BODY", $sformatf("After Finish item Serial transaction: Rx0_p=%b (%0d)",req.Rx0_p, req.Rx0_p), UVM_LOW)
  endtask : body

  // Post body task
  virtual task post_body();
    super.post_body();
  endtask : post_body

endclass : serdes_same_data_for_tx_rx_sequence
