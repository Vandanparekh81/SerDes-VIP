// ------------------------------------------------------------------------ //
// File Name : serdes_parameter_config.sv
// Author Name : Vandan Parekh
// Propetier Name : ASICraft Technologies
// Description : This is serdes_parameter_config class inside this Width 
// parameter is defined which is used in all the components for example in 
// transaction class for declaration of Tx0, Rx0 signals
// ------------------------------------------------------------------------ //

// This parameter is width of parallel signals
parameter WIDTH = 10; 

