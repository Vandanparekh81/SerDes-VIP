// First argument is class name, 
// second arguement is how many times you want to run,
// Third arguement is you want to select random seed(0) or give specific seed(1)
// Fourth arguement is for coverage enable and disable which is disable for only data error injection test
// Fifth arguement is combine all value plus args
serdes_sanity_test 5 0 1 "SCOREBOARD_ENABLE=1 SPEED=1 PARALLEL_TRANSACTION_COUNT=1 SERIAL_TRANSACTION_COUNT=1" 
serdes_sanity_test 1 0 1 "SCOREBOARD_ENABLE=1 SPEED=2 PARALLEL_TRANSACTION_COUNT=1 SERIAL_TRANSACTION_COUNT=1" 
serdes_multiple_transaction_test 1 0 1 "SCOREBOARD_ENABLE=1 SPEED=3 PARALLEL_TRANSACTION_COUNT=5 SERIAL_TRANSACTION_COUNT=2" 
serdes_multiple_transaction_test 1 0 1 "SCOREBOARD_ENABLE=1 SPEED=9 PARALLEL_TRANSACTION_COUNT=8 SERIAL_TRANSACTION_COUNT=5" 
serdes_multiple_transaction_test 1 0 1 "SCOREBOARD_ENABLE=1 SPEED=10 PARALLEL_TRANSACTION_COUNT=9 SERIAL_TRANSACTION_COUNT=6" 
serdes_data_pattern_test 1 0 1 "SCOREBOARD_ENABLE=1 DATA_PATTERN=WALKING_0 SPEED=4 PARALLEL_TRANSACTION_COUNT=20 SERIAL_TRANSACTION_COUNT=20" 
serdes_data_pattern_test 1 0 1 "SCOREBOARD_ENABLE=1 DATA_PATTERN=WALKING_1 SPEED=5 PARALLEL_TRANSACTION_COUNT=10 SERIAL_TRANSACTION_COUNT=15" 
serdes_data_pattern_test 1 0 1 "SCOREBOARD_ENABLE=1 DATA_PATTERN=INCREMENT SPEED=10 PARALLEL_TRANSACTION_COUNT=10 SERIAL_TRANSACTION_COUNT=15" 
serdes_data_pattern_test 1 0 1 "SCOREBOARD_ENABLE=1 DATA_PATTERN=ALTERNATING_5 SPEED=7 PARALLEL_TRANSACTION_COUNT=10 SERIAL_TRANSACTION_COUNT=15" 
serdes_data_pattern_test 5 0 1 "SCOREBOARD_ENABLE=1 DATA_PATTERN=ALTERNATING_A SPEED=8 PARALLEL_TRANSACTION_COUNT=10 SERIAL_TRANSACTION_COUNT=15" 
serdes_data_pattern_test 1 0 1 "SCOREBOARD_ENABLE=1 DATA_PATTERN=ALL_ONE SPEED=9 PARALLEL_TRANSACTION_COUNT=10 SERIAL_TRANSACTION_COUNT=15" 
serdes_data_pattern_test 1 0 1 "SCOREBOARD_ENABLE=1 DATA_PATTERN=ALL_ZERO SPEED=3 PARALLEL_TRANSACTION_COUNT=10 SERIAL_TRANSACTION_COUNT=15" 
serdes_data_pattern_test 1 0 1 "SCOREBOARD_ENABLE=1 DATA_PATTERN=DECREMENT SPEED=2 PARALLEL_TRANSACTION_COUNT=10 SERIAL_TRANSACTION_COUNT=15" 
serdes_data_pattern_test 1 0 1 "SCOREBOARD_ENABLE=1 DATA_PATTERN=RANDOM SPEED=2 PARALLEL_TRANSACTION_COUNT=10 SERIAL_TRANSACTION_COUNT=15" 
serdes_same_data_for_tx_rx_test 1 0 1 "SCOREBOARD_ENABLE=1 SPEED=6 PARALLEL_TRANSACTION_COUNT=20 SERIAL_TRANSACTION_COUNT=20" 
serdes_opposite_data_for_tx_rx_test 1 0 1 "SCOREBOARD_ENABLE=1 SPEED=7 PARALLEL_TRANSACTION_COUNT=18 SERIAL_TRANSACTION_COUNT=18" 
serdes_multiple_transaction_test 1 0 1 "SCOREBOARD_ENABLE=1 SPEED=8 PARALLEL_TRANSACTION_COUNT=5 SERIAL_TRANSACTION_COUNT=2" 
serdes_data_error_injection_test 1 0 0 "SCOREBOARD_ENABLE=1 SPEED=4 PARALLEL_TRANSACTION_COUNT=9 SERIAL_TRANSACTION_COUNT=3" 
