`timescale 1ns/1ps
module sipo_shift_register #(parameter WIDTH=10) 
(
  input logic serial_clk,
  input logic parallel_clk,
  input logic rst,
  input logic Rx0_p, Rx0_n,
  output logic [WIDTH-1 : 0] Rx0
);

  logic [WIDTH-1 : 0] shift_reg;
  logic [WIDTH-1 : 0] parallel_data;
  int sipo_main_count = 0;
  int count = 0;

   always @(posedge serial_clk or posedge rst) begin
    if(rst) begin
      shift_reg <= '0;
      parallel_data <= 0;
      sipo_main_count = 1;
      count = 0;
      `uvm_info("DUT SIPO RESET", $sformatf("RESET CONDITION DISPLAY Serial clock [%0t] Rx0_p = %b | Rx0_p Decimal = %0d |shift_reg = %b | shift_reg in decimal = %0d", $time, Rx0_p, Rx0_p, shift_reg, shift_reg), UVM_LOW)
    end
    else begin
      if(sipo_main_count >= 1) begin
        shift_reg <= {shift_reg[WIDTH-2:0], Rx0_p};
        sipo_main_count++;
        if(count == 0) begin
          if(sipo_main_count == WIDTH+4) begin
            sipo_main_count = 1;
            parallel_data <= shift_reg;
            count++;
          end
        end
        else begin
          if(sipo_main_count == WIDTH+1) begin
            sipo_main_count = 1;
            parallel_data <= shift_reg;
            count++;
          end
        end
      `uvm_info("DUT SIPO", $sformatf("Serial clock [%0t] Rx0_p = %b | Rx0_p Decimal = %0d |shift_reg = %b | shift_reg in decimal = %0d | sipo_main_count = %0d", $time, Rx0_p, Rx0_p, shift_reg, shift_reg, sipo_main_count), UVM_LOW);
      end
      //#1;
    end
  end

  always @(posedge parallel_clk or posedge rst) begin
    if(rst) begin
      sipo_main_count = 1;
      count = 0;
      `uvm_info("DUT SIPO", $sformatf("RESET CONDITION DISPLAY Parallel clock [%0t] Rx0 = %b | Rx0 Decimal = %0d |shift_reg = %b | shift_reg in decimal = %0d", $time, Rx0, Rx0, shift_reg, shift_reg), UVM_LOW)
    end
    else begin 
      //sipo_main_count = 1;
      `uvm_info("DUT SIPO", $sformatf("Parallel clock [%0t] Rx0 = %b | Rx0 Decimal = %0d |shift_reg = %b | shift_reg in decimal = %0d | sipo_main_count = %0d", $time, Rx0, Rx0, shift_reg, shift_reg, sipo_main_count), UVM_LOW)
    end
    end

  assign Rx0 = parallel_data;

   /* always_ff @(posedge serial_clk or posedge rst) begin
    if (rst) begin
      shift_reg <= '0;
      sipo_main_count <= '0;
    end else begin
      shift_reg <= {shift_reg[WIDTH-2:0], Rx0_p}; // shift left
      sipo_main_count <= (sipo_main_count == WIDTH-1) ? 0 : sipo_main_count + 1;
    end
  end

  // Parallel Clock Domain: Capturing 10-bit data after full collection
  always_ff @(posedge parallel_clk or posedge rst) begin
    if (rst) begin
      parallel_data <= '0;
    end else begin
      parallel_data <= shift_reg;
      `uvm_info("DUT SIPO", $sformatf("Parallel clock [%0t] parallel_data = %b | parallel_data Decimal = %0d |shift_reg = %b | shift_reg in decimal = %0d | sipo_main_count = %0d", $time, parallel_data, parallel_data, shift_reg, shift_reg, sipo_main_count), UVM_LOW)
    end
  end

  // Connect to interface output
  assign Rx0 = parallel_data; */

endmodule  



module piso_shift_register #(
    parameter WIDTH = 10 
) (
    input logic serial_clk,
    input logic parallel_clk,
    input logic rst,       
    input logic [WIDTH-1:0] Tx0, 
    output logic Tx0_p, Tx0_n 
);
    logic [WIDTH-1:0] shift_reg;
    int i = 1;
    int count = 0;
    int main_count = 0;


    /* always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            shift_reg <= '0;
        end 
        else if (load) begin
            shift_reg <= Rx0_p;
        end 
        else begin
            shift_reg <= {shift_reg[WIDTH-2:0], 1'b0}; 
        end
    end */

    always @(posedge serial_clk or posedge rst) begin
      if(rst) begin
        Tx0_p <= 0;
        Tx0_n <= 1;
        `uvm_info("DUT PISO RESET CONDITION", $sformatf("RESET CONDITION Serial Clock [%0t] Tx0 = %b | Tx0 Decimal = %0d |Tx0_p = %b | Tx0_n = %0d", $time, Tx0, Tx0, Tx0_p, Tx0_n), UVM_LOW)
      end
      else begin
        if(main_count >= 1) begin 
          Tx0_p <= Tx0[WIDTH-i];
          Tx0_n <= ~Tx0[WIDTH-i];
          `uvm_info("DUT PISO", $sformatf("Serial Clock [%0t] Tx0 = %b | Tx0 Decimal = %0d |Tx0_p = %b | Tx0_n = %0d", $time, Tx0, Tx0, Tx0_p, Tx0_n), UVM_LOW)
          main_count++;
          $display("main_Count = %0d", main_count);
          $display("I = %0d", i);

          if(main_count == WIDTH+1) begin
            main_count = 0;
            i = 1;
          end
          else begin
            i++;
          end
        end

      end
    end

    always @(posedge parallel_clk or posedge rst) begin
      if(rst) begin
        main_count = 0;
      end

      else begin
        main_count = 1;
        //i=0;
      end

    end


endmodule

