class serdes_subscriber extends uvm_subscriber#(serdes_transaction);
   `uvm_component_utils(serdes_subscriber);

  function new (string name, uvm_component parent);
    super.new(name, parent);
  endfunction

  function void build_phase (uvm_phase phase);
    super.build_phase(phase);
  endfunction
