package serdes_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  `include "../seq_lib/serdes_transaction.sv"
  `include "../seq_lib/serdes_sequence.sv"
  `include "serdes_agent_config.sv"
  `include "../test/serdes_test_config.sv"
  `include "../seq_lib/serdes_sequencer.sv"
  `include "serdes_driver.sv"
  `include "serdes_monitor.sv"
  `include "serdes_scoreboard.sv"
  `include "serdes_agent.sv"
  `include "serdes_env.sv"
  `include "../test/serdes_test.sv"
endpackage
import uvm_pkg::*;
`include "uvm_macros.svh"
`include "../../tb_top/serdes_top_tb.sv"
`include "serdes_interface.sv"
`include "../../sve/serdes_dut.sv"
